.TITLE Ex4_1

*****************************
**     Library setting     **
*****************************
.protect
* .include 'Convolution_SYN_new.sp'
.include '7nm_TT.pm'
.include 'asap7sc7p5t_SIMPLE_RVT.sp'
.include 'asap7sc7p5t_SEQ_RVT.sp'
.include 'asap7sc7p5t_OA_RVT.sp'
.include 'asap7sc7p5t_INVBUF_RVT.sp'
.include 'asap7sc7p5t_AO_RVT.sp'
.unprotect

.VEC "Pattern_Convolution.vec"

* .global VDD VSS
Vvdd VDD GND supply
Vvss VSS GND 0

.param supply = 0.75v
* .param total_worktime = 42n


.SUBCKT Convolution VSS VDD  IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Port10
* BUFx10_ASAP7_75t_R VSS VDD A Y
Xbuffer_IFM_03  VSS VDD IFM_0[3] IFM0[3] BUFx10_ASAP7_75t_R
Xbuffer_IFM_02  VSS VDD IFM_0[2] IFM0[2] BUFx10_ASAP7_75t_R
Xbuffer_IFM_01  VSS VDD IFM_0[1] IFM0[1] BUFx10_ASAP7_75t_R
Xbuffer_IFM_00  VSS VDD IFM_0[0] IFM0[0] BUFx10_ASAP7_75t_R

Xbuffer_IFM_13  VSS VDD IFM_1[3] IFM1[3] BUFx10_ASAP7_75t_R
Xbuffer_IFM_12  VSS VDD IFM_1[2] IFM1[2] BUFx10_ASAP7_75t_R
Xbuffer_IFM_11  VSS VDD IFM_1[1] IFM1[1] BUFx10_ASAP7_75t_R
Xbuffer_IFM_10  VSS VDD IFM_1[0] IFM1[0] BUFx10_ASAP7_75t_R

Xbuffer_IFM_23  VSS VDD IFM_2[3] IFM2[3] BUFx10_ASAP7_75t_R
Xbuffer_IFM_22  VSS VDD IFM_2[2] IFM2[2] BUFx10_ASAP7_75t_R
Xbuffer_IFM_21  VSS VDD IFM_2[1] IFM2[1] BUFx10_ASAP7_75t_R
Xbuffer_IFM_20  VSS VDD IFM_2[0] IFM2[0] BUFx10_ASAP7_75t_R

Xbuffer_IFM_33  VSS VDD IFM_3[3] IFM3[3] BUFx10_ASAP7_75t_R
Xbuffer_IFM_32  VSS VDD IFM_3[2] IFM3[2] BUFx10_ASAP7_75t_R
Xbuffer_IFM_31  VSS VDD IFM_3[1] IFM3[1] BUFx10_ASAP7_75t_R
Xbuffer_IFM_30  VSS VDD IFM_3[0] IFM3[0] BUFx10_ASAP7_75t_R

**************************************************
Xbuffer_INW_03  VSS VDD INW_0[3] INW0[3] BUFx10_ASAP7_75t_R
Xbuffer_INW_02  VSS VDD INW_0[2] INW0[2] BUFx10_ASAP7_75t_R
Xbuffer_INW_01  VSS VDD INW_0[1] INW0[1] BUFx10_ASAP7_75t_R
Xbuffer_INW_00  VSS VDD INW_0[0] INW0[0] BUFx10_ASAP7_75t_R

Xbuffer_INW_13  VSS VDD INW_1[3] INW1[3] BUFx10_ASAP7_75t_R
Xbuffer_INW_12  VSS VDD INW_1[2] INW1[2] BUFx10_ASAP7_75t_R
Xbuffer_INW_11  VSS VDD INW_1[1] INW1[1] BUFx10_ASAP7_75t_R
Xbuffer_INW_10  VSS VDD INW_1[0] INW1[0] BUFx10_ASAP7_75t_R

Xbuffer_INW_23  VSS VDD INW_2[3] INW2[3] BUFx10_ASAP7_75t_R
Xbuffer_INW_22  VSS VDD INW_2[2] INW2[2] BUFx10_ASAP7_75t_R
Xbuffer_INW_21  VSS VDD INW_2[1] INW2[1] BUFx10_ASAP7_75t_R
Xbuffer_INW_20  VSS VDD INW_2[0] INW2[0] BUFx10_ASAP7_75t_R

Xbuffer_INW_33  VSS VDD INW_3[3] INW3[3] BUFx10_ASAP7_75t_R
Xbuffer_INW_32  VSS VDD INW_3[2] INW3[2] BUFx10_ASAP7_75t_R
Xbuffer_INW_31  VSS VDD INW_3[1] INW3[1] BUFx10_ASAP7_75t_R
Xbuffer_INW_30  VSS VDD INW_3[0] INW3[0] BUFx10_ASAP7_75t_R

Xmult_18 VSS VDD  IFM0[3] IFM0[2] IFM0[1] IFM0[0] INW0[3] INW0[2] INW0[1] INW0[0] N07 N06 N05 N04 N03 N02 N01 N00 Convolution_DW_mult_uns_3
Xmult_18_2 VSS VDD  IFM1[3] IFM1[2] IFM1[1] IFM1[0] INW1[3] INW1[2] INW1[1] INW1[0] N015 N014 N013 N012 N011 N010 N09 N08 Convolution_DW_mult_uns_2
Xmult_18_3 VSS VDD  IFM2[3] IFM2[2] IFM2[1] IFM2[0] INW2[3] INW2[2] INW2[1] INW2[0] N032 N031 N030 N029 N028 N027 N026 N025 Convolution_DW_mult_uns_1
Xmult_18_4 VSS VDD  IFM3[3] IFM3[2] IFM3[1] IFM3[0] INW3[3] INW3[2] INW3[1] INW3[0] N050 N049 N048 N047 N046 N045 N044 N043 Convolution_DW_mult_uns_0
Xadd_1_root_add_0_root_add_18_3 VSS VDD  N042 N042 N015 N014 N013 N012 N011 N010 N09 N08 N042 N042 N050 N049 N048 N047 N046 N045 N044 N043 N042 SYNOPSYS_UNCONNECTED_1 n9 n8 n7 n6 n5 n4 n3 n2 n1 Convolution_DW01_add_2
Xadd_2_root_add_0_root_add_18_3 VSS VDD  N042 N042 N07 N06 N05 N04 N03 N02 N01 N00 N042 N042 N032 N031 N030 N029 N028 N027 N026 N025 N042 SYNOPSYS_UNCONNECTED_2 N041 N040 N039 N038 N037 N036 N035 N034 N033 Convolution_DW01_add_1
Xadd_0_root_add_0_root_add_18_3 VSS VDD  N042 N041 N040 N039 N038 N037 N036 N035 N034 N033 N042 n9 n8 n7 n6 n5 n4 n3 n2 n1 N042 Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Convolution_DW01_add_0
XU1 VSS VDD  N042 TIELOx1_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW01_add_0 VSS VDD  A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0]
XU1_8 VSS VDD  A[8] B[8] n3 n10 n11 FAx1_ASAP7_75t_R
XU1_7 VSS VDD  A[7] B[7] n4 n12 n13 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n5 n14 n15 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n6 n16 n17 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n7 n18 n19 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n8 n20 n21 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n9 n22 n23 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n24 n25 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n12 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n14 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n16 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n18 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n20 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n22 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n24 n9 INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[9] INVx1_ASAP7_75t_R
XU11 VSS VDD  n11 SUM[8] INVx1_ASAP7_75t_R
XU12 VSS VDD  n13 SUM[7] INVx1_ASAP7_75t_R
XU13 VSS VDD  n15 SUM[6] INVx1_ASAP7_75t_R
XU14 VSS VDD  n17 SUM[5] INVx1_ASAP7_75t_R
XU15 VSS VDD  n19 SUM[4] INVx1_ASAP7_75t_R
XU16 VSS VDD  n21 SUM[3] INVx1_ASAP7_75t_R
XU17 VSS VDD  n23 SUM[2] INVx1_ASAP7_75t_R
XU18 VSS VDD  n25 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW01_add_1 VSS VDD  A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0]
XU1_7 VSS VDD  A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n2 n21 n22 FAx1_ASAP7_75t_R
XU1 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU2 VSS VDD  A[0] B[0] n2 AND2x2_ASAP7_75t_R
XU3 VSS VDD  n11 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n13 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n15 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n17 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n19 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n21 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  n12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  n14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  n16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  n18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW01_add_2 VSS VDD  A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] B[9] B[8] B[7] B[6] B[5] B[4] B[3] B[2] B[1] B[0] CI SUM[9] SUM[8] SUM[7] SUM[6] SUM[5] SUM[4] SUM[3] SUM[2] SUM[1] SUM[0]
XU1_7 VSS VDD  A[7] B[7] n3 n9 n10 FAx1_ASAP7_75t_R
XU1_6 VSS VDD  A[6] B[6] n4 n11 n12 FAx1_ASAP7_75t_R
XU1_5 VSS VDD  A[5] B[5] n5 n13 n14 FAx1_ASAP7_75t_R
XU1_4 VSS VDD  A[4] B[4] n6 n15 n16 FAx1_ASAP7_75t_R
XU1_3 VSS VDD  A[3] B[3] n7 n17 n18 FAx1_ASAP7_75t_R
XU1_2 VSS VDD  A[2] B[2] n8 n19 n20 FAx1_ASAP7_75t_R
XU1_1 VSS VDD  A[1] B[1] n1 n21 n22 FAx1_ASAP7_75t_R
XU1 VSS VDD  A[0] B[0] n1 AND2x2_ASAP7_75t_R
XU2 VSS VDD  B[0] A[0] SUM[0] XOR2xp5_ASAP7_75t_R
XU3 VSS VDD  n11 n3 INVx1_ASAP7_75t_R
XU4 VSS VDD  n13 n4 INVx1_ASAP7_75t_R
XU5 VSS VDD  n15 n5 INVx1_ASAP7_75t_R
XU6 VSS VDD  n17 n6 INVx1_ASAP7_75t_R
XU7 VSS VDD  n19 n7 INVx1_ASAP7_75t_R
XU8 VSS VDD  n21 n8 INVx1_ASAP7_75t_R
XU9 VSS VDD  n9 SUM[8] INVx1_ASAP7_75t_R
XU10 VSS VDD  n10 SUM[7] INVx1_ASAP7_75t_R
XU11 VSS VDD  n12 SUM[6] INVx1_ASAP7_75t_R
XU12 VSS VDD  n14 SUM[5] INVx1_ASAP7_75t_R
XU13 VSS VDD  n16 SUM[4] INVx1_ASAP7_75t_R
XU14 VSS VDD  n18 SUM[3] INVx1_ASAP7_75t_R
XU15 VSS VDD  n20 SUM[2] INVx1_ASAP7_75t_R
XU16 VSS VDD  n22 SUM[1] INVx1_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_0 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_1 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_2 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS


.SUBCKT Convolution_DW_mult_uns_3 VSS VDD  a[3] a[2] a[1] a[0] b[3] b[2] b[1] b[0] product[7] product[6] product[5] product[4] product[3] product[2] product[1] product[0]
XU32 VSS VDD  n41 n44 n31 n25 n26 FAx1_ASAP7_75t_R
XU35 VSS VDD  n36 n45 n32 n29 n30 FAx1_ASAP7_75t_R
XU39 VSS VDD  n49 n52 n38 n34 n35 FAx1_ASAP7_75t_R
XU70 VSS VDD  a[2] n83 INVx1_ASAP7_75t_R
XU71 VSS VDD  n35 n84 INVx1_ASAP7_75t_R
XU72 VSS VDD  a[0] n85 INVx1_ASAP7_75t_R
XU73 VSS VDD  b[3] n86 INVx1_ASAP7_75t_R
XU74 VSS VDD  b[0] n87 INVx1_ASAP7_75t_R
XU75 VSS VDD  n88 n89 product[7] NAND2xp33_ASAP7_75t_R
XU76 VSS VDD  n90 n91 n89 NAND2xp33_ASAP7_75t_R
XU77 VSS VDD  n92 n25 n88 OR2x2_ASAP7_75t_R
XU78 VSS VDD  n91 n90 product[6] XOR2xp5_ASAP7_75t_R
XU79 VSS VDD  n92 n25 n90 XOR2xp5_ASAP7_75t_R
XU80 VSS VDD  b[3] a[3] n92 NAND2xp33_ASAP7_75t_R
XU81 VSS VDD  n93 n94 n91 NAND2xp33_ASAP7_75t_R
XU82 VSS VDD  n95 n96 n94 NAND2xp33_ASAP7_75t_R
XU83 VSS VDD  n26 n29 n93 OR2x2_ASAP7_75t_R
XU84 VSS VDD  n96 n95 product[5] XOR2xp5_ASAP7_75t_R
XU85 VSS VDD  n26 n29 n95 XOR2xp5_ASAP7_75t_R
XU86 VSS VDD  n97 n98 n96 NAND2xp33_ASAP7_75t_R
XU87 VSS VDD  n99 n100 n98 NAND2xp33_ASAP7_75t_R
XU88 VSS VDD  n30 n34 n97 OR2x2_ASAP7_75t_R
XU89 VSS VDD  n100 n99 product[4] XOR2xp5_ASAP7_75t_R
XU90 VSS VDD  n30 n34 n99 XOR2xp5_ASAP7_75t_R
XU91 VSS VDD  n101 n102 n100 NAND2xp33_ASAP7_75t_R
XU92 VSS VDD  n103 n104 n102 NAND2xp33_ASAP7_75t_R
XU93 VSS VDD  n105 n84 n101 NAND2xp33_ASAP7_75t_R
XU94 VSS VDD  n104 n103 product[3] XOR2xp5_ASAP7_75t_R
XU95 VSS VDD  n35 n105 n103 XNOR2xp5_ASAP7_75t_R
XU96 VSS VDD  n106 n107 n105 XOR2xp5_ASAP7_75t_R
XU97 VSS VDD  n108 n109 n104 NAND2xp33_ASAP7_75t_R
XU98 VSS VDD  n110 n111 n109 NAND2xp33_ASAP7_75t_R
XU99 VSS VDD  n112 n113 n108 NAND2xp33_ASAP7_75t_R
XU100 VSS VDD  n110 n111 product[2] XOR2xp5_ASAP7_75t_R
XU101 VSS VDD  n112 n113 n111 XOR2xp5_ASAP7_75t_R
XU102 VSS VDD  n114 n115 n113 XOR2xp5_ASAP7_75t_R
XU103 VSS VDD  n83 n87 n112 NOR2xp33_ASAP7_75t_R
XU104 VSS VDD  n116 n117 n110 NOR2xp33_ASAP7_75t_R
XU105 VSS VDD  n116 n117 product[1] XOR2xp5_ASAP7_75t_R
XU106 VSS VDD  b[1] a[0] n117 NAND2xp33_ASAP7_75t_R
XU107 VSS VDD  b[0] a[1] n116 NAND2xp33_ASAP7_75t_R
XU108 VSS VDD  n87 n85 product[0] NOR2xp33_ASAP7_75t_R
XU109 VSS VDD  n85 n86 n52 NOR2xp33_ASAP7_75t_R
XU110 VSS VDD  a[1] b[2] n49 AND2x2_ASAP7_75t_R
XU111 VSS VDD  a[2] b[2] n45 AND2x2_ASAP7_75t_R
XU112 VSS VDD  n83 n86 n44 NOR2xp33_ASAP7_75t_R
XU113 VSS VDD  b[2] a[3] n41 AND2x2_ASAP7_75t_R
XU114 VSS VDD  n115 n114 n38 NOR2xp33_ASAP7_75t_R
XU115 VSS VDD  b[1] a[1] n114 NAND2xp33_ASAP7_75t_R
XU116 VSS VDD  b[2] a[0] n115 NAND2xp33_ASAP7_75t_R
XU117 VSS VDD  n107 n106 n36 NOR2xp33_ASAP7_75t_R
XU118 VSS VDD  a[3] b[0] n106 NAND2xp33_ASAP7_75t_R
XU119 VSS VDD  a[2] b[1] n107 NAND2xp33_ASAP7_75t_R
XU120 VSS VDD  n118 n119 n32 XOR2xp5_ASAP7_75t_R
XU121 VSS VDD  n118 n119 n31 NOR2xp33_ASAP7_75t_R
XU122 VSS VDD  a[3] b[1] n119 NAND2xp33_ASAP7_75t_R
XU123 VSS VDD  b[3] a[1] n118 NAND2xp33_ASAP7_75t_R
.ENDS

XConvolution VSS VDD IFM_0[3] IFM_0[2] IFM_0[1] IFM_0[0] IFM_1[3] IFM_1[2] IFM_1[1] IFM_1[0] IFM_2[3] IFM_2[2] IFM_2[1] IFM_2[0] IFM_3[3] IFM_3[2] IFM_3[1] IFM_3[0] INW_0[3] INW_0[2] INW_0[1] INW_0[0] INW_1[3] INW_1[2] INW_1[1] INW_1[0] INW_2[3] INW_2[2] INW_2[1] INW_2[0] INW_3[3] INW_3[2] INW_3[1] INW_3[0] Output[9] Output[8] Output[7] Output[6] Output[5] Output[4] Output[3] Output[2] Output[1] Output[0] Port10 Convolution

Cload0 Output[0] VSS 5f
Cload1 Output[1] VSS 5f
Cload2 Output[2] VSS 5f
Cload3 Output[3] VSS 5f
Cload4 Output[4] VSS 5f
Cload5 Output[5] VSS 5f
Cload6 Output[6] VSS 5f
Cload7 Output[7] VSS 5f
Cload8 Output[8] VSS 5f
Cload9 Output[9] VSS 5f


// measurement
.tran 0.1ps 42ns

.measure TRAN Tp1 TRIG V(INW_3[2]) VAL='supply/2'  FALL=1 TARG V(Output[8]) VAL='supply/2'  RISE=1
.measure TRAN Tp2 TRIG V(INW_3[2]) VAL='supply/2'  FALL=2 TARG V(Output[8]) VAL='supply/2'  RISE=2
.measure TRAN Tp3 TRIG V(INW_3[2]) VAL='supply/2'  FALL=3 TARG V(Output[8]) VAL='supply/2'  RISE=3
.measure TRAN Tp4 TRIG V(INW_3[2]) VAL='supply/2'  FALL=4 TARG V(Output[8]) VAL='supply/2'  RISE=4
.measure TRAN Tp5 TRIG V(INW_3[2]) VAL='supply/2'  FALL=5 TARG V(Output[8]) VAL='supply/2'  RISE=5
.measure TRAN Tp6 TRIG V(INW_3[2]) VAL='supply/2'  FALL=6 TARG V(Output[8]) VAL='supply/2'  RISE=6
.measure TRAN Tp7 TRIG V(INW_3[2]) VAL='supply/2'  FALL=7 TARG V(Output[8]) VAL='supply/2'  RISE=7
.measure TRAN Tp8 TRIG V(INW_3[2]) VAL='supply/2'  FALL=8 TARG V(Output[8]) VAL='supply/2'  RISE=8
.measure TRAN Tp9 TRIG V(INW_3[2]) VAL='supply/2'  FALL=9 TARG V(Output[8]) VAL='supply/2'  RISE=9
.measure TRAN Tp10 TRIG V(INW_3[2]) VAL='supply/2'  FALL=10 TARG V(Output[8]) VAL='supply/2'  RISE=10

.measure TRAN Tp11 TRIG V(INW_3[2]) VAL='supply/2'  FALL=11 TARG V(Output[8]) VAL='supply/2'  RISE=11
.measure TRAN Tp12 TRIG V(INW_3[2]) VAL='supply/2'  FALL=12 TARG V(Output[8]) VAL='supply/2'  RISE=12
.measure TRAN Tp13 TRIG V(INW_3[2]) VAL='supply/2'  FALL=13 TARG V(Output[8]) VAL='supply/2'  RISE=13
.measure TRAN Tp14 TRIG V(INW_3[2]) VAL='supply/2'  FALL=14 TARG V(Output[8]) VAL='supply/2'  RISE=14
.measure TRAN Tp15 TRIG V(INW_3[2]) VAL='supply/2'  FALL=15 TARG V(Output[8]) VAL='supply/2'  RISE=15
.measure TRAN Tp16 TRIG V(INW_3[2]) VAL='supply/2'  FALL=16 TARG V(Output[8]) VAL='supply/2'  RISE=17
.measure TRAN Tp17 TRIG V(INW_3[2]) VAL='supply/2'  FALL=17 TARG V(Output[8]) VAL='supply/2'  RISE=18
.measure TRAN Tp18 TRIG V(INW_3[2]) VAL='supply/2'  FALL=18 TARG V(Output[8]) VAL='supply/2'  RISE=19
.measure TRAN Tp19 TRIG V(INW_3[2]) VAL='supply/2'  FALL=19 TARG V(Output[8]) VAL='supply/2'  RISE=20
.measure TRAN Tp20 TRIG V(INW_3[2]) VAL='supply/2'  FALL=20 TARG V(Output[8]) VAL='supply/2'  RISE=21

.measure TRAN average_power avg Power

*****************************
**    Simulator setting    **
*****************************
.op
.option post 
.option probe			*with I/V in .lis
.probe v(*) i(*) 
.option captab			*with cap value in .lis
.TEMP 25


.end